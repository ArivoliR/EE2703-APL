.circuit
V1 1 GND dc 5
R1 1 2 0     # Zero resistance, should be treated as a wire
R2 2 GND 1000
.end

