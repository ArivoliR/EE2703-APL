# Test circuit for negative resistance
.circuit
V1 1 GND dc 5
R1 1 2 1000
R2 2 GND -10   #Negative resistance
.end
